.SUBCKT DFFHQx1 CLK D Q VDD VSS
MM3 pu1 D VDD VNW pmos_lvt l=20n nfin=2
MM1 MH clkb pu1 VNW pmos_lvt l=20n nfin=2
MM5 pd1 D VSS VPW nmos_lvt l=20n nfin=2
MM4 MH clkn pd1 VPW nmos_lvt l=20n nfin=2
MM9 MH clkb pd3 VPW nmos_lvt l=20n nfin=2
MM10 MH clkn pd2 VNW pmos_lvt l=20n nfin=2
MM7 MS MH VDD VNW pmos_lvt l=20n nfin=2
MM6 MS MH VSS VPW nmos_lvt l=20n nfin=2
MM8 pd3 MS VSS VPW nmos_lvt l=20n nfin=2
MM11 pd2 MS VDD VNW pmos_lvt l=20n nfin=2
MM13 MS clkn SH VNW pmos_lvt l=20n nfin=2
MM12 MS clkb SH VPW nmos_lvt l=20n nfin=2
MM20 clkn CLK VSS VPW nmos_lvt l=20n nfin=2
MM23 CLKB clkn VSS VPW nmos_lvt l=20n nfin=2
MM21 clkn CLK VDD VNW pmos_lvt l=20n nfin=2
MM22 CLKB clkn VDD VNW pmos_lvt l=20n nfin=2
MM17 SH clkn pd5 VPW nmos_lvt l=20n nfin=2
MM18 SH clkb pd4 VNW pmos_lvt l=20n nfin=2
MM15 SS SH VDD VNW pmos_lvt l=20n nfin=2
MM14 SS SH VSS VPW nmos_lvt l=20n nfin=2
MM16 pd5 SS VSS VPW nmos_lvt l=20n nfin=2
MM19 pd4 SS VDD VNW pmos_lvt l=20n nfin=2
MM25 Q SS VDD VNW pmos_lvt l=20n nfin=2
MM24 Q SS VSS VPW nmos_lvt l=20n nfin=2
.ENDS


.SUBCKT DFFARHQx1 CLK D RESETN Q VDD VSS
MM21 clkn CLK VDD VNW pmos_lvt l=20n nfin=2
MM22 clkb clkn VDD VNW pmos_lvt l=20n nfin=2
MM20 clkn CLK VSS VPW nmos_lvt l=20n nfin=2
MM23 clkb clkn VSS VPW nmos_lvt l=20n nfin=2
MM1 MH clkb pu1 VNW pmos_lvt l=20n nfin=2
MM3 pu1 D VDD VNW pmos_lvt l=20n nfin=2
MM4 MH clkn pd1 VPW nmos_lvt l=20n nfin=2
MM5 pd1 D VSS VPW nmos_lvt l=20n nfin=2
MM6 VDD MH MS VNW pmos_lvt l=20n nfin=2
MM10 MH clkn net53 VNW pmos_lvt l=20n nfin=2
MM8 VDD MS net53 VNW pmos_lvt l=20n nfin=2
MM11 VDD RESETN net53 VNW pmos_lvt l=20n nfin=2
MM0 net050 RESETN net10 VPW nmos_lvt l=20n nfin=2
MM9 MH clkb net10 VPW nmos_lvt l=20n nfin=2
MM2 VSS MS net050 VPW nmos_lvt l=20n nfin=2
MM46 VSS MH MS VPW nmos_lvt l=20n nfin=2
MM13 MS clkn SH VNW pmos_lvt l=20n nfin=2
MM12 MS clkb SH VPW nmos_lvt l=20n nfin=2
MM24 Q SS VSS VPW nmos_lvt l=20n nfin=2
MM15 net047 RESETN SS VPW nmos_lvt l=20n nfin=2
MM27 VSS SH net047 VPW nmos_lvt l=20n nfin=2
MM18 VSS SS net049 VPW nmos_lvt l=20n nfin=2
MM28 SH clkn net049 VPW nmos_lvt l=20n nfin=2
MM26 VDD RESETN SS VNW pmos_lvt l=20n nfin=2
MM29 SH clkb net030 VNW pmos_lvt l=20n nfin=2
MM25 Q SS VDD VNW pmos_lvt l=20n nfin=2
MM17 VDD SS net030 VNW pmos_lvt l=20n nfin=2
MM19 VDD SH SS VNW pmos_lvt l=20n nfin=2
.ENDS
