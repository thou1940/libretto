.SUBCKT BUFx2 A VDD VPW Y
MM3 Y AN VSS VPW nmos_lvt l=20n nfin=4
MM2 AN A VSS VPW nmos_lvt l=20n nfin=2
MM0 Y AN VDD VNW pmos_lvt l=20n nfin=4
MM1 AN A VDD VNW pmos_lvt l=20n nfin=2
.ENDS


.SUBCKT BUFx3 A VDD VPW Y
MM1 Y AN VDD VNW pmos_lvt l=20n nfin=6
MM0 AN A VDD VNW pmos_lvt l=20n nfin=2
MM2 AN A VSS VPW nmos_lvt l=20n nfin=2
MM3 Y AN VSS VPW nmos_lvt l=20n nfin=6
.ENDS


.SUBCKT BUFx4 A VDD VPW Y
MM1 Y AN VDD VNW pmos_lvt l=20n nfin=8
MM0 AN A VDD VNW pmos_lvt l=20n nfin=2
MM2 AN A VSS VPW nmos_lvt l=20n nfin=2
MM3 Y AN VSS VPW nmos_lvt l=20n nfin=8
.ENDS



.SUBCKT BUFx5 A VDD VPW Y
MM1 Y AN VDD VNW pmos_lvt l=20n nfin=10
MM0 AN A VDD VNW pmos_lvt l=20n nfin=2
MM3 Y AN VSS VPW nmos_lvt l=20n nfin=10
MM2 AN A VSS VPW nmos_lvt l=20n nfin=2
.ENDS


.SUBCKT BUFx6q A VDD VPW Y
MM1 Y AN VDD VNW pmos_lvt l=20n nfin=12
MM0 AN A VDD VNW pmos_lvt l=20n nfin=4
MM3 Y AN VSS VPW nmos_lvt l=20n nfin=12
MM2 AN A VSS VPW nmos_lvt l=20n nfin=4
.ENDS


.SUBCKT BUFx8 A VDD VPW Y
MM0 AN A VDD VNW pmos_lvt l=20n nfin=4
MM1 Y AN VDD VNW pmos_lvt l=20n nfin=16
MM2 AN A VSS VPW nmos_lvt l=20n nfin=4
MM3 Y AN VSS VPW nmos_lvt l=20n nfin=16
.ENDS





