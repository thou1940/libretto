.SUBCKT DFFHQx1 CLK D Q VDD VSS
MM3 pu1 D VDD VDD pmos_lvt l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt l=20n nfin=2
MM4 MH clkn pd1 VSS nmos_lvt l=20n nfin=2
MM9 MH clkb pd3 VSS nmos_lvt l=20n nfin=2
MM10 MH clkn pd2 VDD pmos_lvt l=20n nfin=2
MM7 MS MH VDD VDD pmos_lvt l=20n nfin=2
MM6 MS MH VSS VSS nmos_lvt l=20n nfin=2
MM8 pd3 MS VSS VSS nmos_lvt l=20n nfin=2
MM11 pd2 MS VDD VDD pmos_lvt l=20n nfin=2
MM13 MS clkn SH VDD pmos_lvt l=20n nfin=2
MM12 MS clkb SH VSS nmos_lvt l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt l=20n nfin=2
MM23 CLKB clkn VSS VSS nmos_lvt l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt l=20n nfin=2
MM22 CLKB clkn VDD VDD pmos_lvt l=20n nfin=2
MM17 SH clkn pd5 VSS nmos_lvt l=20n nfin=2
MM18 SH clkb pd4 VDD pmos_lvt l=20n nfin=2
MM15 SS SH VDD VDD pmos_lvt l=20n nfin=2
MM14 SS SH VSS VSS nmos_lvt l=20n nfin=2
MM16 pd5 SS VSS VSS nmos_lvt l=20n nfin=2
MM19 pd4 SS VDD VDD pmos_lvt l=20n nfin=2
MM25 Q SS VDD VDD pmos_lvt l=20n nfin=2
MM24 Q SS VSS VSS nmos_lvt l=20n nfin=2
.ENDS



.SUBCKT DFFARHQx1 CLK D RESETN Q VDD VSS
MM21 clkn CLK VDD VDD pmos_lvt l=20n nfin=2
MM22 clkb clkn VDD VDD pmos_lvt l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt l=20n nfin=2
MM23 clkb clkn VSS VSS nmos_lvt l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt l=20n nfin=2
MM3 pu1 D VDD VDD pmos_lvt l=20n nfin=2
MM4 MH clkn pd1 VSS nmos_lvt l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt l=20n nfin=2
MM6 VDD MH MS VDD pmos_lvt l=20n nfin=2
MM10 MH clkn net53 VDD pmos_lvt l=20n nfin=2
MM8 VDD MS net53 VDD pmos_lvt l=20n nfin=2
MM11 VDD RESETN net53 VDD pmos_lvt l=20n nfin=2
MM0 net050 RESETN net10 VSS nmos_lvt l=20n nfin=2
MM9 MH clkb net10 VSS nmos_lvt l=20n nfin=2
MM2 VSS MS net050 VSS nmos_lvt l=20n nfin=2
MM46 VSS MH MS VSS nmos_lvt l=20n nfin=2
MM13 MS clkn SH VDD pmos_lvt l=20n nfin=2
MM12 MS clkb SH VSS nmos_lvt l=20n nfin=2
MM24 Q SS VSS VSS nmos_lvt l=20n nfin=2
MM15 net047 RESETN SS VSS nmos_lvt l=20n nfin=2
MM27 VSS SH net047 VSS nmos_lvt l=20n nfin=2
MM18 VSS SS net049 VSS nmos_lvt l=20n nfin=2
MM28 SH clkn net049 VSS nmos_lvt l=20n nfin=2
MM26 VDD RESETN SS VDD pmos_lvt l=20n nfin=2
MM29 SH clkb net030 VDD pmos_lvt l=20n nfin=2
MM25 Q SS VDD VDD pmos_lvt l=20n nfin=2
MM17 VDD SS net030 VDD pmos_lvt l=20n nfin=2
MM19 VDD SH SS VDD pmos_lvt l=20n nfin=2
.ENDS
