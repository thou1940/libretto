.SUBCKT XOR2x1 A B VDD VSS Y
MM4 VDD A net019 VDD pmos_lvt l=20n nfin=2
MM5 VDD B net019 VDD pmos_lvt l=20n nfin=2
MM6 net019 net036 Y VDD pmos_lvt l=20n nfin=2
MM2 net048 B net036 VDD pmos_lvt l=20n nfin=2
MM3 VDD A net048 VDD pmos_lvt l=20n nfin=2
MM11 VSS A net047 VSS nmos_lvt l=20n nfin=2
MM10 net047 B Y VSS nmos_lvt l=20n nfin=2
MM9 VSS net036 Y VSS nmos_lvt l=20n nfin=2
MM0 VSS A net036 VSS nmos_lvt l=20n nfin=2
MM1 VSS B net036 VSS nmos_lvt l=20n nfin=2
.ENDS


.SUBCKT XOR2x2 A B VDD VSS Y
MM6 xor net067 net071 VSS nmos_lvt l=20n nfin=2
MM2 net067 B net079 VSS nmos_lvt l=20n nfin=2
MM13 VSS xor Y VSS nmos_lvt l=20n nfin=4
MM5 net071 B VSS VSS nmos_lvt l=20n nfin=2
MM3 net079 A VSS VSS nmos_lvt l=20n nfin=2
MM4 net071 A VSS VSS nmos_lvt l=20n nfin=2
MM10 xor B net078 VDD pmos_lvt l=20n nfin=2
MM1 net067 B VDD VDD pmos_lvt l=20n nfin=2
MM12 VDD xor Y VDD pmos_lvt l=20n nfin=4
MM0 net067 A VDD VDD pmos_lvt l=20n nfin=2
MM9 xor net067 VDD VDD pmos_lvt l=20n nfin=2
MM11 net078 A VDD VDD pmos_lvt l=20n nfin=2
.ENDS