.model nmos_lvt nmos (BULKMOD=1 CDSC=0.0242792648477108 CDSCD=0.00392734735055704 CFD=0 CFS=0 CGDL=2.46057180997666e-10 CGDO=0 CGEOMOD=0 CGSL=2.46057180997666e-10 CGSO=0 CIT=0 CJSWGD=5.57527110441952e-11 CJSWGS=5.57527110441952e-11 CKAPPAD=1 CKAPPAS=1 DELVFBACC=0.343773452656344 DSUB=0.938843990618648 DVT0=1e-05 DVT1=0.6 EOT=7.42868560178388e-10 EOTACC=4.71671117014025e-10 ETA0=0.660104661399005 ETAMOB=2 EU=1.44812928246679 GEOMOD=1 HFIN=6e-09 Imin=1e-15 KSATIV=10 L=1.9e-08 MEXP=2.8151407047218 NBODY=3e+24 NFIN=1 NSD=8e+26 NSDE=3e+25 PCLM=0.005 PCLMG=0 PHIG=4.24998827791051 PTWG=0 QMFACTOR=1 QMFACTORCV=1 QMTCENCVA=0 RDSW=22.5584908190333 RGEOMOD=0 TFIN=5.7e-08 TYPE=1 U0=0.0301122423249245 UA=0.616262044625125 VFBSD=0 VFBSDCV=-0.4 VSAT=52245.0479995332 VSAT1=74377.1574945721 level=110)