.SUBCKT AND2x2 A B VNW VSS Y
MM4 Y net10 VDD VNW pmos_lvt l=20n nfin=4
MM1 net10 B VDD VNW pmos_lvt l=20n nfin=2
MM0 net10 A VDD VNW pmos_lvt l=20n nfin=2
MM5 Y net10 VSS VPW nmos_lvt l=20n nfin=4
MM3 net20 A VSS VPW nmos_lvt l=20n nfin=2
MM2 net10 B net20 VPW nmos_lvt l=20n nfin=2
.ENDS


.SUBCKT AND2x4 A B VNW VSS Y
MM4 Y net9 VDD VNW pmos_lvt l=20n nfin=8
MM1 net9 B VDD VNW pmos_lvt l=20n nfin=4
MM0 net9 A VDD VNW pmos_lvt l=20n nfin=4
MM5 Y net9 VSS VPW nmos_lvt l=20n nfin=8
MM3 net19 A VSS VPW nmos_lvt l=20n nfin=4
MM2 net9 B net19 VPW nmos_lvt l=20n nfin=4
.ENDS


.SUBCKT AND2x6 A B VNW VSS Y
MM4 Y net9 VDD VNW pmos_lvt l=20n nfin=12
MM1 net9 B VDD VNW pmos_lvt l=20n nfin=4
MM0 net9 A VDD VNW pmos_lvt l=20n nfin=4
MM5 Y net9 VSS VPW nmos_lvt l=20n nfin=12
MM3 net19 A VSS VPW nmos_lvt l=20n nfin=4
MM2 net9 B net19 VPW nmos_lvt l=20n nfin=4
.ENDS
