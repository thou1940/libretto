.model pmos_lvt pmos (BULKMOD=1 CDSC=0.0298779937685466 CDSCD=0.00592672124113853 CFD=0 CFS=0 CGDL=2.32284344700851e-10 CGDO=0 CGEOMOD=0 CGSL=2.32284344700851e-10 CGSO=0 CIT=0 CJSWGD=4.2579335429074e-11 CJSWGS=4.2579335429074e-11 CKAPPAD=0.707838632342404 CKAPPAS=0.707838632342404 DELVFBACC=0.493819530768007 DSUB=0.855490406783821 DVT0=1e-05 DVT1=0.6 EOT=4.96372131536353e-10 EOTACC=4.58991464641434e-10 ETA0=0.684038031113596 ETAMOB=2 EU=3.07677593816472 GEOMOD=1 HFIN=6e-09 Imin=1e-15 KSATIV=10 L=1.9e-08 MEXP=2.87983831737946 NBODY=3e+24 NFIN=1 NSD=8e+26 NSDE=3e+25 PCLM=0.005 PCLMG=0 PHIG=4.9237703205239 PTWG=0 QMFACTOR=1 QMFACTORCV=1 QMTCENCVA=0 RDSW=1 RGEOMOD=0 TFIN=5.7e-08 TYPE=0 U0=0.0247936000247227 UA=1.40724669571314 VFBSD=0 VFBSDCV=-0.363815960677205 VSAT=80555.5289404872 VSAT1=48818.3387050927 level=110)