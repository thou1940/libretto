.SUBCKT AOI21x1 A1 A2 B VDD VSS Y
MM4 Y B VSS VSS nmos_lvt l=20n nfin=2
MM3 Y A1 net29 VSS nmos_lvt l=20n nfin=2
MM2 net29 A2 VSS VSS nmos_lvt l=20n nfin=2
MM5 net18 A2 VDD VDD pmos_lvt l=20n nfin=2
MM0 Y B net18 VDD pmos_lvt l=20n nfin=2
MM1 net18 A1 VDD VDD pmos_lvt l=20n nfin=2
.ENDS


.SUBCKT AOI21x2 A1 A2 B VDD VSS Y
MM4 Y B VSS VSS nmos_lvt l=20n nfin=4
MM3 Y A1 net29 VSS nmos_lvt l=20n nfin=4
MM2 net29 A2 VSS VSS nmos_lvt l=20n nfin=4
MM5 net18 A2 VDD VDD pmos_lvt l=20n nfin=4
MM0 Y B net18 VDD pmos_lvt l=20n nfin=4
MM1 net18 A1 VDD VDD pmos_lvt l=20n nfin=4
.ENDS

.SUBCKT AOI22xp5 A1 A2 B1 B2 VDD VSS Y
MM5 Y A2 net13 VDD pmos_lvt l=20n nfin=2
MM4 Y A1 net13 VDD pmos_lvt l=20n nfin=2
MM3 net13 B2 VDD VDD pmos_lvt l=20n nfin=2
MM2 net13 B1 VDD VDD pmos_lvt l=20n nfin=2
MM9 net29 B1 VSS VSS nmos_lvt l=20n nfin=2
MM8 net30 A1 VSS VSS nmos_lvt l=20n nfin=2
MM7 Y B2 net29 VSS nmos_lvt l=20n nfin=2
MM6 Y A2 net30 VSS nmos_lvt l=20n nfin=2
.ENDS